package states_pkg;
  typedef enum {INIT,DECODE,IDLE} fmstate_e;
  bit running = 1;
endpackage

